* EESchema Netlist Version 1.1 (Spice format) creation date: 12/15/2014 4:07:39 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  2 3 VPLOT8		
v1  1 0 SINE		
U1  1 VPLOT8_1		
R1  2 3 10k		
D4  0 2 1n4007		
D3  3 0 1n4007		
D2  1 2 1n4007		
D1  3 1 1n4007		

.end
